package core_pkg;

endpackage : mini_dbg_pkg
